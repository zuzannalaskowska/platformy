���      �sklearn.linear_model._logistic��LogisticRegression���)��}�(�penalty��l2��dual���tol�G?6��C-�C�G?�      �fit_intercept���intercept_scaling�K�class_weight�N�random_state�N�solver��lbfgs��max_iter�M��multi_class��auto��verbose�K �
warm_start���n_jobs�N�l1_ratio�N�n_features_in_�K	�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����u1�����R�(K�|�NNNJ����J����K t�b�C �t�b�n_iter_�hhK ��h ��R�(KK��h%�i4�����R�(K�<�NNNJ����J����K t�b�CZ  �t�b�coef_�hhK ��h ��R�(KKK	��h%�f8�����R�(Kh5NNNJ����J����K t�b�CH�ǚ^�B?��mB��?�p����S7�){)"�з4�!�/��r�\?�(@����?uy��g�����~4c�9?�t�b�
intercept_�hhK ��h ��R�(KK��h@�C~H���ڢ��t�b�_sklearn_version��0.24.2�ub.